package shared_pkg;

logic error_cnt;
logic correct_cnt;
bit test_finished;
event sample_event;

endpackage : shared_pkg